`timescale 1ns / 1ps

module gremlin_rom
    (
        input  wire        clk,
        input  wire [2:0] addr1,
        input wire [4:0] addr2,            // {char_code[6:0], char_line[3:0]}
        output wire  [15:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [15:0] data;

    // body
assign char_line_pixels = data;


    always @*
        case (addr2 + (addr1*32))
            //code 000
            8'b000_00000: data = 16'b0000001111000000; //      ****
            8'b000_00001: data = 16'b0000111111110000; //    ********
            8'b000_00010: data = 16'b0001111111111000; //   **********
            8'b000_00011: data = 16'b0001111111111000; //   **********
            8'b000_00100: data = 16'b0001111111111000; //   **********
            8'b000_00101: data = 16'b0000111111110000; //    ********
            8'b000_00110: data = 16'b0000000111000000; //       ***
            8'b000_00111: data = 16'b0000000111000000; //       ***
            8'b000_01000: data = 16'b0000111111110000; //    ********
            8'b000_01001: data = 16'b0011111111111100; //  ************
            8'b000_01010: data = 16'b0111111111111100; // *************
            8'b000_01011: data = 16'b1111111111111100; //**************
            8'b000_01100: data = 16'b1101111111111110; //** ************
            8'b000_01101: data = 16'b1001111111111110; //*  ************
            8'b000_01110: data = 16'b0001111111111110; //   ************
            8'b000_01111: data = 16'b0001111111111010; //   ********** *
            8'b000_10000: data = 16'b0001111111111000; //   **********
            8'b000_10001: data = 16'b0001111111111000; //   **********
            8'b000_10010: data = 16'b0001111111111000; //   **********
            8'b000_10011: data = 16'b0001111111111000; //   **********
            8'b000_10100: data = 16'b0001111111111000; //   **********
            8'b000_10101: data = 16'b0001111111111000; //   **********
            8'b000_10110: data = 16'b0001111111111000; //   **********
            8'b000_10111: data = 16'b0001111111111000; //   **********
            8'b000_11000: data = 16'b0000111001110000; //    ***  ***
            8'b000_11001: data = 16'b0000111000111000; //    ***   ***
            8'b000_11010: data = 16'b0000111000011100; //    ***    ***
            8'b000_11011: data = 16'b0000011000001110; //     **     ***
            8'b000_11100: data = 16'b0000011000000111; //     **      ***
            8'b000_11101: data = 16'b0000011000001111; //     **     ****
            8'b000_11110: data = 16'b0000111000001110; //    ***     ***
            8'b000_11111: data = 16'b0000111000000000; //    ***
            //code 001
            8'b001_00000: data = 16'b0000001111000000; //      ****
            8'b001_00001: data = 16'b0000111111110000; //    ********
            8'b001_00010: data = 16'b0001111111111000; //   **********
            8'b001_00011: data = 16'b0001111111111000; //   **********
            8'b001_00100: data = 16'b0001111111111000; //   **********
            8'b001_00101: data = 16'b0000111111110000; //    ********
            8'b001_00110: data = 16'b0000000111000000; //       ***
            8'b001_00111: data = 16'b0000000111000000; //       ***
            8'b001_01000: data = 16'b0000111111110000; //    ********
            8'b001_01001: data = 16'b1111111111111100; //**************
            8'b001_01010: data = 16'b1111111111111110; //***************
            8'b001_01011: data = 16'b1111111111111111; //****************
            8'b001_01100: data = 16'b0001111111111011; //   ********** **
            8'b001_01101: data = 16'b0001111111111001; //   **********  *
            8'b001_01110: data = 16'b0001111111111000; //   **********
            8'b001_01111: data = 16'b0001111111111000; //   **********   
            8'b001_10000: data = 16'b0001111111111000; //   **********
            8'b001_10001: data = 16'b0001111111111000; //   **********
            8'b001_10010: data = 16'b0001111111111000; //   **********
            8'b001_10011: data = 16'b0001111111111000; //   **********
            8'b001_10100: data = 16'b0001111111111000; //   **********
            8'b001_10101: data = 16'b0001111111111000; //   **********
            8'b001_10110: data = 16'b0001111111111000; //   **********
            8'b001_10111: data = 16'b0001111111111000; //   **********
            8'b001_11000: data = 16'b0000111001110000; //    ***  ***   
            8'b001_11001: data = 16'b0001110001110000; //   ***   ***    
            8'b001_11010: data = 16'b0011100001110000; //  ***    ***
            8'b001_11011: data = 16'b0111000000111000; // ***      ***
            8'b001_11100: data = 16'b0111000000011100; // ***       ***
            8'b001_11101: data = 16'b0110000000001100; // **         **     
            8'b001_11110: data = 16'b1110000000011100; //***        ***
            8'b001_11111: data = 16'b1110000000011100; //***        ***
            //code x02
            8'b001_00000: data = 16'b0000000000000000; //  
            8'b001_00001: data = 16'b0000000000000000; //
            8'b001_00010: data = 16'b0000000000000000; //
            8'b001_00011: data = 16'b0000000000000000; //
            8'b001_00100: data = 16'b0000000000000000; //
            8'b001_00101: data = 16'b0000000000000000; //
            8'b001_00110: data = 16'b0000000000000000; //
            8'b001_00111: data = 16'b0000000000000000; //
            8'b001_01000: data = 16'b0000000000000000; //
            8'b001_01001: data = 16'b0000000000000000; //
            8'b001_01010: data = 16'b0000000000000000; //
            8'b001_01011: data = 16'b0000000000000000; //
            8'b001_01100: data = 16'b0000000000000000; //
            8'b001_01101: data = 16'b0000000000000000; //
            8'b001_01110: data = 16'b0000000000000000; //
            8'b001_01111: data = 16'b0000000000000000; //   
            8'b001_10000: data = 16'b0000000000000000; //    
            8'b001_10001: data = 16'b0000000000000000; //    
            8'b001_10010: data = 16'b0000000000000000; //    
            8'b001_10011: data = 16'b0000000000000000; //    
            8'b001_10100: data = 16'b0000000000000000; //     
            8'b001_10101: data = 16'b0000000000000000; //    
            8'b001_10110: data = 16'b0000000000000000; //     
            8'b001_10111: data = 16'b0000000000000000; //      
            8'b001_11000: data = 16'b0000000000000000; //   
            8'b001_11001: data = 16'b0000000000000000; //    
            8'b001_11010: data = 16'b0000000000000000; //     
            8'b001_11011: data = 16'b0000000000000000; //     
            8'b001_11100: data = 16'b0000000000000000; //      
            8'b001_11101: data = 16'b0000000000000000; //     
            8'b001_11110: data = 16'b0000000000000000; //     
            8'b001_11111: data = 16'b0000000000000000; //
            //code x03
            8'b000_00000: data = 16'b0000001111000000; //      ****
            8'b000_00001: data = 16'b0000001111000000; //      ****
            8'b000_00010: data = 16'b0000001111000000; //      ****
            8'b000_00011: data = 16'b0000001111000000; //      ****
            8'b000_00100: data = 16'b0000001111000000; //      ****
            8'b000_00101: data = 16'b0000001111000000; //      ****
            8'b000_00110: data = 16'b1111111111111111; //****************
            8'b000_00111: data = 16'b1111111111111111; //****************
            8'b000_01000: data = 16'b1111111111111111; //****************
            8'b000_01001: data = 16'b1111111111111111; //****************
            8'b000_01010: data = 16'b0000001111000000; //      ****
            8'b000_01011: data = 16'b0000001111000000; //      ****
            8'b000_01100: data = 16'b0000001111000000; //      ****
            8'b000_01101: data = 16'b0000001111000000; //      ****
            8'b000_01110: data = 16'b0000001111000000; //      ****
            8'b000_01111: data = 16'b0000001111000000; //      ****
            8'b000_10000: data = 16'b0000001111000000; //      ****
            8'b000_10001: data = 16'b0000001111000000; //      ****
            8'b000_10010: data = 16'b0000001111000000; //      ****
            8'b000_10011: data = 16'b0000001111000000; //      ****
            8'b000_10100: data = 16'b0000001111000000; //      ****
            8'b000_10101: data = 16'b0000001111000000; //      ****
            8'b000_10110: data = 16'b0000001111000000; //      ****
            8'b000_10111: data = 16'b0000001111000000; //      ****
            8'b000_11000: data = 16'b0000001111000000; //      ****
            8'b000_11001: data = 16'b0000001111000000; //      ****
            8'b000_11010: data = 16'b0000001111000000; //      ****
            8'b000_11011: data = 16'b0000001111000000; //      ****
            8'b000_11100: data = 16'b0000001111000000; //      ****
            8'b000_11101: data = 16'b0000001111000000; //      ****
            8'b000_11110: data = 16'b1111111111111111; //****************
            8'b000_11111: data = 16'b1111111111111111; //****************
            //code x04
        endcase

endmodule
