`timescale 1ns / 1ps

module gremlin_rom
    (
        input wire addr1,
        input wire [4:0] addr2,            // {char_code[6:0], char_line[3:0]}
        output wire  [15:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [15:0] data;

    // body
assign char_line_pixels = data;


    always @*
        case (addr2 + (addr1*32))
            //code 000
            6'b0_00000: data = 16'b0000001111000000; //      ****
            6'b0_00001: data = 16'b0000111111110000; //    ********
            6'b0_00010: data = 16'b0001111111111000; //   **********
            6'b0_00011: data = 16'b0001111111111000; //   **********
            6'b0_00100: data = 16'b0001111111111000; //   **********
            6'b0_00101: data = 16'b0000111111110000; //    ********
            6'b0_00110: data = 16'b0000000111000000; //       ***
            6'b0_00111: data = 16'b0000000111000000; //       ***
            6'b0_01000: data = 16'b0000111111110000; //    ********
            6'b0_01001: data = 16'b0011111111111100; //  ************
            6'b0_01010: data = 16'b0111111111111100; // *************
            6'b0_01011: data = 16'b1111111111111100; //**************
            6'b0_01100: data = 16'b1101111111111110; //** ************
            6'b0_01101: data = 16'b1001111111111110; //*  ************
            6'b0_01110: data = 16'b0001111111111110; //   ************
            6'b0_01111: data = 16'b0001111111111010; //   ********** *
            6'b0_10000: data = 16'b0001111111111000; //   **********
            6'b0_10001: data = 16'b0001111111111000; //   **********
            6'b0_10010: data = 16'b0001111111111000; //   **********
            6'b0_10011: data = 16'b0001111111111000; //   **********
            6'b0_10100: data = 16'b0001111111111000; //   **********
            6'b0_10101: data = 16'b0001111111111000; //   **********
            6'b0_10110: data = 16'b0001111111111000; //   **********
            6'b0_10111: data = 16'b0001111111111000; //   **********
            6'b0_11000: data = 16'b0000111001110000; //    ***  ***
            6'b0_11001: data = 16'b0000111000111000; //    ***   ***
            6'b0_11010: data = 16'b0000111000011100; //    ***    ***
            6'b0_11011: data = 16'b0000011000001110; //     **     ***
            6'b0_11100: data = 16'b0000011000000111; //     **      ***
            6'b0_11101: data = 16'b0000011000001111; //     **     ****
            6'b0_11110: data = 16'b0000111000001110; //    ***     ***
            6'b0_11111: data = 16'b0000111000000000; //    ***
            //code 001
            6'b1_00000: data = 16'b0000001111000000; //      ****
            6'b1_00001: data = 16'b0000111111110000; //    ********
            6'b1_00010: data = 16'b0001111111111000; //   **********
            6'b1_00011: data = 16'b0001111111111000; //   **********
            6'b1_00100: data = 16'b0001111111111000; //   **********
            6'b1_00101: data = 16'b0000111111110000; //    ********
            6'b1_00110: data = 16'b0000000111000000; //       ***
            6'b1_00111: data = 16'b0000000111000000; //       ***
            6'b1_01000: data = 16'b0000111111110000; //    ********
            6'b1_01001: data = 16'b1111111111111100; //**************
            6'b1_01010: data = 16'b1111111111111110; //***************
            6'b1_01011: data = 16'b1111111111111111; //****************
            6'b1_01100: data = 16'b0001111111111011; //   ********** **
            6'b1_01101: data = 16'b0001111111111001; //   **********  *
            6'b1_01110: data = 16'b0001111111111000; //   **********
            6'b1_01111: data = 16'b0001111111111000; //   **********   
            6'b1_10000: data = 16'b0001111111111000; //   **********
            6'b1_10001: data = 16'b0001111111111000; //   **********
            6'b1_10010: data = 16'b0001111111111000; //   **********
            6'b1_10011: data = 16'b0001111111111000; //   **********
            6'b1_10100: data = 16'b0001111111111000; //   **********
            6'b1_10101: data = 16'b0001111111111000; //   **********
            6'b1_10110: data = 16'b0001111111111000; //   **********
            6'b1_10111: data = 16'b0001111111111000; //   **********
            6'b1_11000: data = 16'b0000111001110000; //    ***  ***   
            6'b1_11001: data = 16'b0001110001110000; //   ***   ***    
            6'b1_11010: data = 16'b0011100001110000; //  ***    ***
            6'b1_11011: data = 16'b0111000000111000; // ***      ***
            6'b1_11100: data = 16'b0111000000011100; // ***       ***
            6'b1_11101: data = 16'b0110000000001100; // **         **     
            6'b1_11110: data = 16'b1110000000011100; //***        ***
            6'b1_11111: data = 16'b1110000000011100; //***        ***

        endcase

endmodule
